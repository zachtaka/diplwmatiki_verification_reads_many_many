/** 
 * @info Master NI
 * 
 * @author VLSI Lab, EE dept., Democritus University of Thrace
 * 
 * @brief The Master NI contains:
 *        (a) Buffers for AXI AW, W, B and R channels (removed appropriately if Write or Read channels are not present)
 *        (b) Request path, which is followed by transactions, upont exiting the NoC (@see axi_master_ni_req_path),
 *            to feed the external Slave's AW, W and AR channels.
 *        (c) Response path, which is followed by response transactions generated by the external Slave at the B and R channels
 *            (@see axi_slave_ni_resp_path)
 *
 * @param SLAVE_ID specifies the ID of the External Slave, attached to the Master NI
 * @param TIDS_M specifies the number of AXI Transaction IDs at the External Master Side
 * @param ADDRESS_WIDTH specifies the address filed width of the transactions (AxADDR)
 * @param DATA_LANES specifies the number of byte lanes of the Write Data channel (W)
 * @param USER_WIDTH specifies the width of the US field of the AXI channels
 * @param EXT_MASTERS specifies the number of the system's External Masters
 * @param EXT_SLAVES specifies the number of External AXI Slave
 * @param HAS_WRITE specifies if the NI serves Write Requests (simplifies unit if it doesn't)
 * @param HAS_READ specifies if the NI serves Read Requests (simplifies unit if it doesn't)
 * @param MAX_LINK_WIDTH_REQ specifies the maximum tolerated link width of the NoC request path (@see axi_master_ni_req_path)
 * @param MAX_LINK_WIDTH_RESP specifies the maximum tolerated link width of the NoC response path (@see axi_resp_packetizer)
 * @param AW_FIFO_DEPTH specifies the buffer slots of the AW channel output FIFO buffer
 * @param W_FIFO_DEPTH specifies the buffer slots of the W channel output FIFO buffer
 * @param AR_FIFO_DEPTH specifies the buffer slots of the AR channel output FIFO buffer
 * @param B_FIFO_DEPTH specifies the buffer slots of the B channel input FIFO buffer
 * @param R_FIFO_DEPTH specifies the buffer slots of the R channel input FIFO buffer
 * @param FLIT_WIDTH_REQ_C specifies the width of the request flit.
 * @param FLIT_WIDTH_RESP_C specifies the width of the response.
 * @param NI_NOC_FC_SND specifies buffering and flow control (@see flow_control_sender) of the NI->NoC link (response path)
 * @param NOC_NI_FC_RCV specifies buffering and flow control (@see flow_control_receiver) of the NoC->NI link (request path)
 */

import axi4_duth_noc_pkg::*;
import axi4_duth_noc_ni_pkg::*;


module axi_master_ni
  #(parameter int SLAVE_ID                              = 0,
    parameter int TIDS_M                                = 16,
    parameter int ADDRESS_WIDTH                         = 32,
    parameter int DATA_LANES                            = 4,
    parameter int USER_WIDTH                            = 2,
    parameter int EXT_MASTERS                           = 4,
    parameter int EXT_SLAVES                            = 2,
    parameter logic HAS_WRITE                           = 1'b1,
    parameter logic HAS_READ                            = 1'b1,
    parameter int MAX_LINK_WIDTH_REQ                    = 128,
    parameter int MAX_LINK_WIDTH_RESP                   = 128,
    parameter int AW_FIFO_DEPTH                         = 2,
    parameter int W_FIFO_DEPTH                          = 2,
    parameter int AR_FIFO_DEPTH                         = 2,
    parameter int B_FIFO_DEPTH                          = 2,
    parameter int R_FIFO_DEPTH                          = 2,
    // Flit widths passed here to avoid recaclulation
    parameter int FLIT_WIDTH_REQ_C                      = 128,
    parameter int FLIT_WIDTH_RESP_C                     = 128,
    parameter link_fc_params_snd_type NI_NOC_FC_SND     = RTR_CREDITS_3_FC_SND,
    parameter link_fc_params_rcv_type NOC_NI_FC_RCV     = RTR_CREDITS_3_FC_RCV,
    parameter logic ASSERT_RV               = 1'b0)
   (input logic clk,
    input logic rst,
    ///   NoC Side   ///
    // NoC -> Req flits
    input logic[FLIT_WIDTH_REQ_C-1 : 0] req_flit_from_noc,
    input logic req_valid_from_noc,
    output logic req_ready_to_noc,
    // NoC <- Resp Flits
    output logic[FLIT_WIDTH_RESP_C-1 : 0] resp_flit_to_noc,
    output logic resp_valid_to_noc,
    input logic resp_ready_from_noc,
    ///   Slave Side   ///
    // Write Address
    output logic[log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + ADDRESS_WIDTH + USER_WIDTH + AXI_W_AWR_STD_FIELDS-1 : 0] aw_chan,
    output logic aw_valid,
    input logic aw_ready,
    // Write Data
    output logic[log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + 9*DATA_LANES + USER_WIDTH + AXI_SPECS_WIDTH_LAST-1 : 0] w_chan,
    output logic w_valid,
    input logic w_ready,
    // Read Address
    output logic[log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + ADDRESS_WIDTH + USER_WIDTH + AXI_W_AWR_STD_FIELDS-1 : 0] ar_chan,
    output logic ar_valid,
    input logic ar_ready,
    // Write Response
    input logic[log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + USER_WIDTH + AXI_SPECS_WIDTH_RESP-1 : 0] b_chan,
    input logic b_valid,
    output logic b_ready,
    // Read Data
    input logic[log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + 8*DATA_LANES + USER_WIDTH + AXI_SPECS_WIDTH_RESP + AXI_SPECS_WIDTH_LAST-1 : 0] r_chan,
    input logic r_valid,
    output logic r_ready);


// pragma synthesis_off
// pragma translate_off
initial begin
    $display("FIFOs @ Master NI %0d (AW, W, B, AR, R: %0d %0d %0d %0d %0d)", SLAVE_ID,  AW_FIFO_DEPTH, W_FIFO_DEPTH, B_FIFO_DEPTH, AR_FIFO_DEPTH, R_FIFO_DEPTH);
end
// pragma synthesis_on
// pragma translate_on
    
// Slave Side Channel Widths (outgoing)
localparam AXI_W_AWR_S = log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + ADDRESS_WIDTH + USER_WIDTH + AXI_W_AWR_STD_FIELDS;
localparam AXI_W_W_S   = log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + 9*DATA_LANES + USER_WIDTH + AXI_SPECS_WIDTH_LAST;
localparam AXI_W_B_S   = log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + USER_WIDTH + AXI_SPECS_WIDTH_RESP;
localparam AXI_W_R_S   = log2c_1if1(TIDS_M) + $clog2(EXT_MASTERS) + 8*DATA_LANES + USER_WIDTH + AXI_SPECS_WIDTH_RESP + AXI_SPECS_WIDTH_LAST;

// Ready/Valid monitoring
// AW
rv_handshake_checker
        #(  .DATA_WIDTH (AXI_W_AWR_S),
            .ASSERT_EN  (ASSERT_RV))
    rv_mon_aw
        (   .clk    (clk),
            .rst    (rst),
            .data   (aw_chan),
            .valid  (aw_valid),
            .ready  (aw_ready));
// W
rv_handshake_checker
        #(  .DATA_WIDTH (AXI_W_W_S),
            .ASSERT_EN  (ASSERT_RV))
    rv_mon_w
        (   .clk    (clk),
            .rst    (rst),
            .data   (w_chan),
            .valid  (w_valid),
            .ready  (w_ready));
// AR
rv_handshake_checker
        #(  .DATA_WIDTH (AXI_W_AWR_S),
            .ASSERT_EN  (ASSERT_RV))
    rv_mon_ar
        (   .clk    (clk),
            .rst    (rst),
            .data   (ar_chan),
            .valid  (ar_valid),
            .ready  (ar_ready));
// B
rv_handshake_checker
        #(  .DATA_WIDTH (AXI_W_B_S),
            .ASSERT_EN  (ASSERT_RV))
    rv_mon_b
        (   .clk    (clk),
            .rst    (rst),
            .data   (b_chan),
            .valid  (b_valid),
            .ready  (b_ready));
// R
rv_handshake_checker
        #(  .DATA_WIDTH (AXI_W_R_S),
            .ASSERT_EN  (ASSERT_RV))
    rv_mon_r
        (   .clk    (clk),
            .rst    (rst),
            .data   (r_chan),
            .valid  (r_valid),
            .ready  (r_ready));

// NoC Channel Input Queue
logic[FLIT_WIDTH_REQ_C-1 : 0] noc_req_fifo_data;
logic noc_req_fifo_valid, noc_req_fifo_ready;
    
// AXI Output Queues
// AW
logic[AXI_W_AWR_S-1 : 0] aw_fifo_data;
logic aw_fifo_ready, aw_fifo_valid;
// W
logic[AXI_W_W_S-1 : 0] w_fifo_data;
logic w_fifo_ready, w_fifo_valid;
/// AR
logic[AXI_W_AWR_S-1 : 0] ar_fifo_data;
logic ar_fifo_ready, ar_fifo_valid;
    
// AXI Input Queues
// B
logic[AXI_W_B_S-1 : 0] b_fifo_data;
logic b_fifo_ready, b_fifo_valid;
// R
logic[AXI_W_R_S-1 : 0] r_fifo_data;
logic r_fifo_ready, r_fifo_valid;
    
// NoC Channel Output Queue
logic[FLIT_WIDTH_RESP_C-1 : 0] noc_resp_fifo_data;
logic noc_resp_fifo_ready, noc_resp_fifo_valid;

// Work-around for tool unsupporting on-the-fly enum assignment
localparam link_fc_params_snd_type AW_FC_SND_PARAMS = '{FC_TYPE:FLOW_CONTROL_ELASTIC, PUSH_CHECK_READY: 1'b1, CR_MAX_CREDITS:3, CR_REG_DATA:1'b0, CR_REG_CR_UPD:1'b0, CR_USE_INCR:1'b0, RV_BUFF_DEPTH:AW_FIFO_DEPTH};
localparam link_fc_params_snd_type W_FC_SND_PARAMS  = '{FC_TYPE:FLOW_CONTROL_ELASTIC, PUSH_CHECK_READY: 1'b1, CR_MAX_CREDITS:3, CR_REG_DATA:1'b0, CR_REG_CR_UPD:1'b0, CR_USE_INCR:1'b0, RV_BUFF_DEPTH:W_FIFO_DEPTH};
localparam link_fc_params_snd_type AR_FC_SND_PARAMS = '{FC_TYPE:FLOW_CONTROL_ELASTIC, PUSH_CHECK_READY: 1'b1, CR_MAX_CREDITS:3, CR_REG_DATA:1'b0, CR_REG_CR_UPD:1'b0, CR_USE_INCR:1'b0, RV_BUFF_DEPTH:AR_FIFO_DEPTH};
localparam link_fc_params_rcv_type B_FC_RCV_PARAMS  = '{FC_TYPE:FLOW_CONTROL_ELASTIC, BUFF_DEPTH:B_FIFO_DEPTH, POP_CHECK_VALID:1'b1, CR_REG_CR_UPD:1'b0, RV_PUSH_CHECK_READY:1'b1};
localparam link_fc_params_rcv_type R_FC_RCV_PARAMS  = '{FC_TYPE:FLOW_CONTROL_ELASTIC, BUFF_DEPTH:R_FIFO_DEPTH, POP_CHECK_VALID:1'b1, CR_REG_CR_UPD:1'b0, RV_PUSH_CHECK_READY:1'b1};

// NoC Input Buffer
flow_control_receiver #(.LINK_WIDTH         (FLIT_WIDTH_REQ_C),
                        .FC_RCV_PARAMS		(NOC_NI_FC_RCV))
inp_buf_noc_req(.clk              (clk),
                .rst              (rst),
                .data_in          (req_flit_from_noc),
                .valid_in         (req_valid_from_noc),
                .back_notify      (req_ready_to_noc),
                .data_out         (noc_req_fifo_data),
                .valid_out        (noc_req_fifo_valid),
                .ready_in         (noc_req_fifo_ready));

// Request NI
axi_master_ni_req_path #(.SLAVE_ID             (SLAVE_ID),
                         .TIDS_M               (TIDS_M),
                         .ADDRESS_WIDTH        (ADDRESS_WIDTH),
                         .DATA_LANES           (DATA_LANES),
                         .USER_WIDTH           (USER_WIDTH),
                         .EXT_MASTERS          (EXT_MASTERS),
                         .EXT_SLAVES           (EXT_SLAVES),
                         .MAX_LINK_WIDTH_REQ   (MAX_LINK_WIDTH_REQ),
                         .FLIT_WIDTH_REQ_C     (FLIT_WIDTH_REQ_C))
noc_to_s_ni(.clk             (clk),
            .rst             (rst),
            .inp_chan        (noc_req_fifo_data),
            .inp_valid       (noc_req_fifo_valid),
            .inp_ready       (noc_req_fifo_ready),
            .aw_chan         (aw_fifo_data),
            .aw_valid        (aw_fifo_valid),
            .aw_ready        (aw_fifo_ready),
            .w_chan          (w_fifo_data),
            .w_valid         (w_fifo_valid),
            .w_ready         (w_fifo_ready),
            .ar_chan         (ar_fifo_data),
            .ar_valid        (ar_fifo_valid),
            .ar_ready        (ar_fifo_ready));
            
            

generate
  // AXI Output Buffering
  if (HAS_WRITE) begin
    if (AW_FIFO_DEPTH > 0) begin: aw_fc
          // AW
          flow_control_sender #(.LINK_WIDTH         (AXI_W_AWR_S),
                                .FC_SND_PARAMS		(AW_FC_SND_PARAMS))
          out_buf_axi_aw(.clk              (clk),
                         .rst              (rst),
                         .data_in          (aw_fifo_data),
                         .valid_in         (aw_fifo_valid),
                         .ready_out        (aw_fifo_ready),
                         .data_out         (aw_chan),
                         .valid_out        (aw_valid),
                         .front_notify     (aw_ready));
    end else begin: aw_dum
        assign aw_chan = aw_fifo_data;
        assign aw_valid = aw_fifo_valid;
        assign aw_fifo_ready = aw_ready;
    end
    
    if (W_FIFO_DEPTH > 0) begin: w_fc
          // W
          flow_control_sender #(.LINK_WIDTH         (AXI_W_W_S),
                                .FC_SND_PARAMS		    (W_FC_SND_PARAMS))
          out_buf_axi_w(.clk              (clk),
                        .rst              (rst),
                        .data_in          (w_fifo_data),
                        .valid_in         (w_fifo_valid),
                        .ready_out        (w_fifo_ready),
                        .data_out         (w_chan),
                        .valid_out        (w_valid),
                        .front_notify     (w_ready));
    end else begin: w_dum
        assign w_chan = w_fifo_data;
        assign w_valid = w_fifo_valid;
        assign w_fifo_ready = w_ready;
    end
  end else begin
    //NOT HAS_WRITE
      assign aw_valid = 0;
      assign aw_fifo_ready = 0;
      assign w_valid  = 0;
      assign w_fifo_ready  = 0;
    end
    
  if (HAS_READ)
    if (AR_FIFO_DEPTH > 0) begin: ar_fc
        // AR
        flow_control_sender #(.LINK_WIDTH         (AXI_W_AWR_S),
                              .FC_SND_PARAMS	  (AR_FC_SND_PARAMS))
        out_buf_axi_ar(.clk              (clk),
                       .rst              (rst),
                       .data_in          (ar_fifo_data),
                       .valid_in         (ar_fifo_valid),
                       .ready_out        (ar_fifo_ready),
                       .data_out         (ar_chan),
                       .valid_out        (ar_valid),
                       .front_notify     (ar_ready));
    end else begin: ar_dum
        assign ar_chan = ar_fifo_data;
        assign ar_valid = ar_fifo_valid;
        assign ar_fifo_ready = ar_ready;
    end
  else begin
    //NOT HAS_READ
      assign ar_valid = 0;
      assign ar_fifo_ready = 0;
    end

        
  // AXI Input Buffering
  if (HAS_WRITE)
    if (B_FIFO_DEPTH > 0) begin: b_fc
        // B
        flow_control_receiver #(.LINK_WIDTH         (AXI_W_B_S),
                                .FC_RCV_PARAMS		 (B_FC_RCV_PARAMS))
        inp_buf_axi_b(.clk              (clk),
                      .rst              (rst),
                      .data_in          (b_chan),
                      .valid_in         (b_valid),
                      .back_notify      (b_ready),
                      .data_out         (b_fifo_data),
                      .valid_out        (b_fifo_valid),
                      .ready_in         (b_fifo_ready));
    end else begin: b_dum
        assign b_fifo_data = b_chan;
        assign b_fifo_valid = b_valid;
        assign b_ready = b_fifo_ready;
    end
  else
    // NOT HAS_WRITE
    begin
      assign b_ready = 0;
      assign b_fifo_valid = 0;
    end
        
  if (HAS_READ)
    if (R_FIFO_DEPTH > 0) begin: r_fc
        // R
        flow_control_receiver #(.LINK_WIDTH         (AXI_W_R_S),
                                .FC_RCV_PARAMS		 (R_FC_RCV_PARAMS))
        inp_buf_axi_r(.clk              (clk),
                      .rst              (rst),
                      .data_in          (r_chan),
                      .valid_in         (r_valid),
                      .back_notify      (r_ready),
                      .data_out         (r_fifo_data),
                      .valid_out        (r_fifo_valid),
                      .ready_in         (r_fifo_ready));
    end else begin: r_dum
        assign r_fifo_data = r_chan;
        assign r_fifo_valid = r_valid;
        assign r_ready = r_fifo_ready;
    end
  else
    // NOT HAS_READ
    begin
      assign r_ready = 0;
      assign r_fifo_valid = 0;
    end

  // Response NI
  axi_master_ni_resp_path #(.SLAVE_ID             (SLAVE_ID), 
                            .TIDS_M               (TIDS_M), 
                            .ADDRESS_WIDTH        (ADDRESS_WIDTH), 
                            .DATA_LANES           (DATA_LANES), 
                            .USER_WIDTH           (USER_WIDTH), 
                            .EXT_MASTERS          (EXT_MASTERS), 
                            .EXT_SLAVES           (EXT_SLAVES),  
                            .HAS_WRITE            (HAS_WRITE), 
                            .HAS_READ             (HAS_READ),
                            .MAX_LINK_WIDTH_RESP  (MAX_LINK_WIDTH_RESP), 
                            .FLIT_WIDTH_C         (FLIT_WIDTH_RESP_C))
  s_to_noc_ni(.clk           (clk), 
              .rst           (rst),
              .b_chan        (b_fifo_data),
              .b_valid       (b_fifo_valid),
              .b_ready       (b_fifo_ready),
              .r_chan        (r_fifo_data),
              .r_valid       (r_fifo_valid),
              .r_ready       (r_fifo_ready),
              .outp_chan     (noc_resp_fifo_data),
              .outp_valid    (noc_resp_fifo_valid),
              .outp_ready    (noc_resp_fifo_ready));
    
  // NoC Output Buffer
  flow_control_sender #(.LINK_WIDTH         (FLIT_WIDTH_RESP_C),
						.FC_SND_PARAMS		(NI_NOC_FC_SND))
  out_buf_noc_resp(.clk              (clk),
                   .rst              (rst),
                   .data_in          (noc_resp_fifo_data),
                   .valid_in         (noc_resp_fifo_valid),
                   .ready_out        (noc_resp_fifo_ready),
                   .data_out         (resp_flit_to_noc),
                   .valid_out        (resp_valid_to_noc),
                   .front_notify     (resp_ready_from_noc));  

endgenerate 
  
endmodule
